magic
tech sky130A
timestamp 1617762838
<< nwell >>
rect 570 -540 1260 -385
rect 1060 -610 1260 -540
<< nmos >>
rect 640 -775 655 -675
rect 705 -775 720 -675
rect 850 -775 865 -675
rect 1020 -775 1035 -675
rect 1085 -775 1100 -675
rect 1260 -775 1275 -675
rect 1325 -775 1340 -675
rect 705 -1025 720 -925
rect 770 -1025 785 -925
rect 835 -1025 850 -925
rect 900 -1025 915 -925
rect 965 -1025 980 -925
rect 1030 -1025 1045 -925
rect 1095 -1025 1110 -925
rect 1160 -1025 1175 -925
<< pmos >>
rect 640 -510 655 -410
rect 705 -510 720 -410
rect 850 -510 865 -410
rect 915 -510 930 -410
rect 1110 -510 1125 -410
rect 1175 -510 1190 -410
<< ndiff >>
rect 590 -690 640 -675
rect 590 -760 605 -690
rect 625 -760 640 -690
rect 590 -775 640 -760
rect 655 -690 705 -675
rect 655 -760 670 -690
rect 690 -760 705 -690
rect 655 -775 705 -760
rect 720 -690 770 -675
rect 720 -760 735 -690
rect 755 -760 770 -690
rect 720 -775 770 -760
rect 800 -690 850 -675
rect 800 -760 815 -690
rect 835 -760 850 -690
rect 800 -775 850 -760
rect 865 -690 915 -675
rect 865 -760 880 -690
rect 900 -760 915 -690
rect 865 -775 915 -760
rect 970 -690 1020 -675
rect 970 -760 985 -690
rect 1005 -760 1020 -690
rect 970 -775 1020 -760
rect 1035 -690 1085 -675
rect 1035 -760 1050 -690
rect 1070 -760 1085 -690
rect 1035 -775 1085 -760
rect 1100 -690 1150 -675
rect 1100 -760 1115 -690
rect 1135 -760 1150 -690
rect 1100 -775 1150 -760
rect 1210 -690 1260 -675
rect 1210 -760 1225 -690
rect 1245 -760 1260 -690
rect 1210 -775 1260 -760
rect 1275 -690 1325 -675
rect 1275 -760 1290 -690
rect 1310 -760 1325 -690
rect 1275 -775 1325 -760
rect 1340 -690 1390 -675
rect 1340 -760 1355 -690
rect 1375 -760 1390 -690
rect 1340 -775 1390 -760
rect 655 -940 705 -925
rect 655 -1010 670 -940
rect 690 -1010 705 -940
rect 655 -1025 705 -1010
rect 720 -940 770 -925
rect 720 -1010 735 -940
rect 755 -1010 770 -940
rect 720 -1025 770 -1010
rect 785 -940 835 -925
rect 785 -1010 800 -940
rect 820 -1010 835 -940
rect 785 -1025 835 -1010
rect 850 -940 900 -925
rect 850 -1010 865 -940
rect 885 -1010 900 -940
rect 850 -1025 900 -1010
rect 915 -940 965 -925
rect 915 -1010 930 -940
rect 950 -1010 965 -940
rect 915 -1025 965 -1010
rect 980 -940 1030 -925
rect 980 -1010 995 -940
rect 1015 -1010 1030 -940
rect 980 -1025 1030 -1010
rect 1045 -940 1095 -925
rect 1045 -1010 1060 -940
rect 1080 -1010 1095 -940
rect 1045 -1025 1095 -1010
rect 1110 -940 1160 -925
rect 1110 -1010 1125 -940
rect 1145 -1010 1160 -940
rect 1110 -1025 1160 -1010
rect 1175 -940 1225 -925
rect 1175 -1010 1190 -940
rect 1210 -1010 1225 -940
rect 1175 -1025 1225 -1010
<< pdiff >>
rect 590 -425 640 -410
rect 590 -495 605 -425
rect 625 -495 640 -425
rect 590 -510 640 -495
rect 655 -425 705 -410
rect 655 -495 670 -425
rect 690 -495 705 -425
rect 655 -510 705 -495
rect 720 -425 770 -410
rect 720 -495 735 -425
rect 755 -495 770 -425
rect 720 -510 770 -495
rect 800 -425 850 -410
rect 800 -495 815 -425
rect 835 -495 850 -425
rect 800 -510 850 -495
rect 865 -425 915 -410
rect 865 -495 880 -425
rect 900 -495 915 -425
rect 865 -510 915 -495
rect 930 -425 980 -410
rect 930 -495 945 -425
rect 965 -495 980 -425
rect 930 -510 980 -495
rect 1060 -425 1110 -410
rect 1060 -495 1075 -425
rect 1095 -495 1110 -425
rect 1060 -510 1110 -495
rect 1125 -425 1175 -410
rect 1125 -495 1140 -425
rect 1160 -495 1175 -425
rect 1125 -510 1175 -495
rect 1190 -425 1240 -410
rect 1190 -495 1205 -425
rect 1225 -495 1240 -425
rect 1190 -510 1240 -495
<< ndiffc >>
rect 605 -760 625 -690
rect 670 -760 690 -690
rect 735 -760 755 -690
rect 815 -760 835 -690
rect 880 -760 900 -690
rect 985 -760 1005 -690
rect 1050 -760 1070 -690
rect 1115 -760 1135 -690
rect 1225 -760 1245 -690
rect 1290 -760 1310 -690
rect 1355 -760 1375 -690
rect 670 -1010 690 -940
rect 735 -1010 755 -940
rect 800 -1010 820 -940
rect 865 -1010 885 -940
rect 930 -1010 950 -940
rect 995 -1010 1015 -940
rect 1060 -1010 1080 -940
rect 1125 -1010 1145 -940
rect 1190 -1010 1210 -940
<< pdiffc >>
rect 605 -495 625 -425
rect 670 -495 690 -425
rect 735 -495 755 -425
rect 815 -495 835 -425
rect 880 -495 900 -425
rect 945 -495 965 -425
rect 1075 -495 1095 -425
rect 1140 -495 1160 -425
rect 1205 -495 1225 -425
<< psubdiff >>
rect 630 -595 730 -580
rect 630 -615 645 -595
rect 715 -615 730 -595
rect 630 -630 730 -615
rect 1195 -820 1295 -805
rect 1195 -840 1210 -820
rect 1280 -840 1295 -820
rect 1195 -855 1295 -840
rect 605 -940 655 -925
rect 605 -1010 620 -940
rect 640 -1010 655 -940
rect 605 -1025 655 -1010
<< nsubdiff >>
rect 1100 -555 1200 -540
rect 1100 -575 1115 -555
rect 1185 -575 1200 -555
rect 1100 -590 1200 -575
<< psubdiffcont >>
rect 645 -615 715 -595
rect 1210 -840 1280 -820
rect 620 -1010 640 -940
<< nsubdiffcont >>
rect 1115 -575 1185 -555
<< poly >>
rect 595 -365 635 -355
rect 595 -385 605 -365
rect 625 -380 635 -365
rect 625 -385 720 -380
rect 595 -395 720 -385
rect 640 -410 655 -395
rect 705 -410 720 -395
rect 850 -410 865 -395
rect 915 -400 1190 -385
rect 915 -410 930 -400
rect 1110 -410 1125 -400
rect 1175 -410 1190 -400
rect 640 -525 655 -510
rect 705 -525 720 -510
rect 850 -525 865 -510
rect 915 -525 930 -510
rect 1110 -525 1125 -510
rect 1175 -525 1190 -510
rect 805 -560 845 -550
rect 805 -580 815 -560
rect 835 -575 845 -560
rect 835 -580 950 -575
rect 805 -590 950 -580
rect 1215 -550 1255 -540
rect 1215 -570 1225 -550
rect 1245 -570 1255 -550
rect 1215 -580 1255 -570
rect 640 -675 655 -660
rect 705 -675 720 -660
rect 850 -675 865 -660
rect 640 -790 655 -775
rect 705 -790 720 -775
rect 850 -790 865 -775
rect 705 -800 910 -790
rect 705 -805 880 -800
rect 870 -820 880 -805
rect 900 -820 910 -800
rect 870 -830 910 -820
rect 935 -855 950 -590
rect 1415 -605 1455 -595
rect 1415 -620 1425 -605
rect 1020 -625 1425 -620
rect 1445 -625 1455 -605
rect 1020 -635 1455 -625
rect 1020 -675 1035 -635
rect 1085 -675 1100 -660
rect 1260 -675 1275 -660
rect 1325 -675 1340 -660
rect 1020 -790 1035 -775
rect 1085 -790 1100 -775
rect 1260 -790 1275 -775
rect 1325 -790 1340 -775
rect 975 -800 1035 -790
rect 975 -820 985 -800
rect 1005 -805 1035 -800
rect 1060 -800 1100 -790
rect 1005 -820 1015 -805
rect 975 -830 1015 -820
rect 1060 -820 1070 -800
rect 1090 -820 1100 -800
rect 1325 -800 1365 -790
rect 1060 -830 1100 -820
rect 1325 -820 1335 -800
rect 1355 -820 1365 -800
rect 1325 -830 1365 -820
rect 900 -870 950 -855
rect 1135 -870 1175 -860
rect 705 -925 720 -910
rect 770 -925 785 -910
rect 835 -925 850 -910
rect 900 -925 915 -870
rect 1135 -890 1145 -870
rect 1165 -890 1175 -870
rect 1135 -900 1175 -890
rect 965 -925 980 -910
rect 1030 -925 1045 -910
rect 1095 -925 1110 -910
rect 1160 -925 1175 -900
rect 705 -1040 720 -1025
rect 770 -1040 785 -1025
rect 835 -1040 850 -1025
rect 900 -1040 915 -1025
rect 965 -1040 980 -1025
rect 1030 -1040 1045 -1025
rect 1095 -1040 1110 -1025
rect 1160 -1040 1175 -1025
rect 705 -1055 1175 -1040
<< polycont >>
rect 605 -385 625 -365
rect 815 -580 835 -560
rect 1225 -570 1245 -550
rect 880 -820 900 -800
rect 1425 -625 1445 -605
rect 985 -820 1005 -800
rect 1070 -820 1090 -800
rect 1335 -820 1355 -800
rect 1145 -890 1165 -870
<< locali >>
rect 595 -365 635 -355
rect 595 -385 605 -365
rect 625 -385 635 -365
rect 595 -395 635 -385
rect 595 -415 615 -395
rect 595 -425 635 -415
rect 595 -495 605 -425
rect 625 -495 635 -425
rect 595 -505 635 -495
rect 660 -425 700 -415
rect 660 -495 670 -425
rect 690 -495 700 -425
rect 660 -505 700 -495
rect 725 -425 765 -415
rect 725 -495 735 -425
rect 755 -495 765 -425
rect 725 -505 765 -495
rect 595 -680 615 -505
rect 635 -595 725 -585
rect 635 -615 645 -595
rect 715 -615 725 -595
rect 635 -625 725 -615
rect 670 -680 690 -625
rect 745 -680 765 -505
rect 805 -425 845 -415
rect 805 -495 815 -425
rect 835 -495 845 -425
rect 805 -505 845 -495
rect 870 -425 910 -415
rect 870 -495 880 -425
rect 900 -495 910 -425
rect 870 -505 910 -495
rect 935 -425 975 -415
rect 935 -495 945 -425
rect 965 -495 975 -425
rect 935 -505 975 -495
rect 805 -550 825 -505
rect 955 -550 975 -505
rect 805 -560 845 -550
rect 805 -580 815 -560
rect 835 -580 845 -560
rect 805 -590 845 -580
rect 890 -570 975 -550
rect 1065 -425 1105 -415
rect 1065 -495 1075 -425
rect 1095 -495 1105 -425
rect 1065 -505 1105 -495
rect 1130 -425 1170 -415
rect 1130 -495 1140 -425
rect 1160 -495 1170 -425
rect 1130 -505 1170 -495
rect 1195 -425 1235 -415
rect 1195 -495 1205 -425
rect 1225 -485 1235 -425
rect 1225 -495 1385 -485
rect 1195 -505 1385 -495
rect 890 -680 910 -570
rect 1065 -595 1085 -505
rect 1140 -545 1160 -505
rect 1105 -555 1195 -545
rect 1105 -575 1115 -555
rect 1185 -575 1195 -555
rect 1105 -585 1195 -575
rect 1215 -550 1255 -540
rect 1215 -570 1225 -550
rect 1245 -570 1255 -550
rect 1215 -580 1255 -570
rect 595 -690 635 -680
rect 595 -760 605 -690
rect 625 -760 635 -690
rect 595 -770 635 -760
rect 660 -690 700 -680
rect 660 -760 670 -690
rect 690 -760 700 -690
rect 660 -770 700 -760
rect 725 -690 765 -680
rect 725 -760 735 -690
rect 755 -760 765 -690
rect 725 -770 765 -760
rect 805 -690 845 -680
rect 805 -760 815 -690
rect 835 -760 845 -690
rect 805 -770 845 -760
rect 870 -690 910 -680
rect 870 -760 880 -690
rect 900 -760 910 -690
rect 870 -770 910 -760
rect 890 -790 910 -770
rect 870 -800 910 -790
rect 870 -820 880 -800
rect 900 -820 910 -800
rect 870 -830 910 -820
rect 975 -615 1085 -595
rect 975 -680 995 -615
rect 1215 -680 1235 -580
rect 1365 -680 1385 -505
rect 1415 -605 1455 -595
rect 1415 -625 1425 -605
rect 1445 -615 1455 -605
rect 1445 -625 1470 -615
rect 1415 -635 1470 -625
rect 975 -690 1015 -680
rect 975 -760 985 -690
rect 1005 -760 1015 -690
rect 975 -770 1015 -760
rect 1040 -690 1080 -680
rect 1040 -760 1050 -690
rect 1070 -760 1080 -690
rect 1040 -770 1080 -760
rect 1105 -690 1145 -680
rect 1105 -760 1115 -690
rect 1135 -750 1145 -690
rect 1215 -690 1255 -680
rect 1215 -750 1225 -690
rect 1135 -760 1225 -750
rect 1245 -760 1255 -690
rect 1105 -770 1255 -760
rect 1280 -690 1320 -680
rect 1280 -760 1290 -690
rect 1310 -760 1320 -690
rect 1280 -770 1320 -760
rect 1345 -690 1385 -680
rect 1345 -760 1355 -690
rect 1375 -760 1385 -690
rect 1345 -770 1385 -760
rect 975 -790 995 -770
rect 1060 -790 1080 -770
rect 975 -800 1015 -790
rect 975 -820 985 -800
rect 1005 -820 1015 -800
rect 975 -830 1015 -820
rect 1060 -800 1100 -790
rect 1060 -820 1070 -800
rect 1090 -820 1100 -800
rect 1280 -810 1300 -770
rect 1345 -790 1365 -770
rect 1060 -830 1100 -820
rect 1200 -820 1300 -810
rect 1200 -840 1210 -820
rect 1280 -840 1300 -820
rect 1325 -800 1365 -790
rect 1325 -820 1335 -800
rect 1355 -810 1365 -800
rect 1355 -820 1470 -810
rect 1325 -830 1470 -820
rect 1200 -850 1300 -840
rect 1135 -870 1175 -860
rect 1135 -880 1145 -870
rect 735 -890 1145 -880
rect 1165 -890 1175 -870
rect 735 -900 1175 -890
rect 735 -930 755 -900
rect 865 -930 885 -900
rect 995 -930 1015 -900
rect 1125 -930 1145 -900
rect 610 -940 700 -930
rect 610 -1010 620 -940
rect 640 -1010 670 -940
rect 690 -1010 700 -940
rect 610 -1020 700 -1010
rect 725 -940 765 -930
rect 725 -1010 735 -940
rect 755 -1010 765 -940
rect 725 -1020 765 -1010
rect 790 -940 830 -930
rect 790 -1010 800 -940
rect 820 -1010 830 -940
rect 790 -1020 830 -1010
rect 855 -940 895 -930
rect 855 -1010 865 -940
rect 885 -1010 895 -940
rect 855 -1020 895 -1010
rect 920 -940 960 -930
rect 920 -1010 930 -940
rect 950 -1010 960 -940
rect 920 -1020 960 -1010
rect 985 -940 1025 -930
rect 985 -1010 995 -940
rect 1015 -1010 1025 -940
rect 985 -1020 1025 -1010
rect 1050 -940 1090 -930
rect 1050 -1010 1060 -940
rect 1080 -1010 1090 -940
rect 1050 -1020 1090 -1010
rect 1115 -940 1155 -930
rect 1115 -1010 1125 -940
rect 1145 -1010 1155 -940
rect 1115 -1020 1155 -1010
rect 1180 -940 1220 -930
rect 1180 -1010 1190 -940
rect 1210 -1010 1220 -940
rect 1180 -1020 1220 -1010
rect 670 -1040 690 -1020
rect 800 -1040 820 -1020
rect 930 -1040 950 -1020
rect 1060 -1040 1080 -1020
rect 1190 -1040 1210 -1020
rect 670 -1060 1210 -1040
<< viali >>
rect 670 -495 690 -425
rect 880 -495 900 -425
rect 1140 -495 1160 -425
rect 1225 -570 1245 -550
rect 670 -760 690 -690
rect 815 -760 835 -690
rect 1050 -760 1070 -690
rect 1290 -760 1310 -690
rect 670 -1010 690 -940
<< metal1 >>
rect 570 -425 1260 -410
rect 570 -495 670 -425
rect 690 -495 880 -425
rect 900 -495 1140 -425
rect 1160 -495 1260 -425
rect 570 -510 1260 -495
rect 1215 -550 1260 -510
rect 1215 -570 1225 -550
rect 1245 -570 1260 -550
rect 1215 -590 1260 -570
rect 575 -690 1400 -675
rect 575 -760 670 -690
rect 690 -760 815 -690
rect 835 -760 1050 -690
rect 1070 -760 1290 -690
rect 1310 -760 1400 -690
rect 575 -775 1400 -760
rect 655 -940 705 -775
rect 655 -1010 670 -940
rect 690 -1010 705 -940
rect 655 -1025 705 -1010
<< labels >>
rlabel metal1 570 -460 570 -460 7 VP
port 7 w
rlabel metal1 575 -730 575 -730 7 VN
port 6 w
rlabel locali 1470 -820 1470 -820 3 VBN
port 4 e
rlabel locali 1470 -625 1470 -625 3 VG
port 3 e
<< end >>
