magic
tech sky130A
timestamp 1617739874
<< error_p >>
rect 2445 -600 2495 -100
rect 3695 -600 3745 -100
<< nmos >>
rect -5 -600 1195 -100
rect 1245 -600 2445 -100
rect 2495 -600 3695 -100
<< ndiff >>
rect -55 -115 -5 -100
rect -55 -585 -40 -115
rect -20 -585 -5 -115
rect -55 -600 -5 -585
rect 1195 -115 1245 -100
rect 1195 -585 1210 -115
rect 1230 -585 1245 -115
rect 1195 -600 1245 -585
rect 2445 -115 2495 -100
rect 2445 -585 2460 -115
rect 2480 -585 2495 -115
rect 2445 -600 2495 -585
rect 3695 -115 3745 -100
rect 3695 -585 3710 -115
rect 3730 -585 3745 -115
rect 3695 -600 3745 -585
<< ndiffc >>
rect -40 -585 -20 -115
rect 1210 -585 1230 -115
rect 2460 -585 2480 -115
rect 3710 -585 3730 -115
<< psubdiff >>
rect -105 -115 -55 -100
rect -105 -585 -90 -115
rect -70 -585 -55 -115
rect -105 -600 -55 -585
<< psubdiffcont >>
rect -90 -585 -70 -115
<< poly >>
rect -55 -55 -15 -45
rect -55 -75 -45 -55
rect -25 -70 -15 -55
rect -25 -75 1195 -70
rect -55 -85 1195 -75
rect -5 -100 1195 -85
rect 1245 -100 2445 -85
rect 2495 -100 3695 -85
rect -5 -615 1195 -600
rect 1245 -615 2445 -600
rect 2495 -615 3695 -600
<< polycont >>
rect -45 -75 -25 -55
<< locali >>
rect -55 -55 -15 -45
rect -55 -75 -45 -55
rect -25 -75 -15 -55
rect -55 -85 -15 -75
rect -50 -105 -30 -85
rect -100 -115 -10 -105
rect -100 -585 -90 -115
rect -70 -585 -40 -115
rect -20 -585 -10 -115
rect -100 -595 -10 -585
rect 1200 -115 1240 -105
rect 1200 -585 1210 -115
rect 1230 -585 1240 -115
rect 1200 -595 1240 -585
rect 2450 -115 2490 -105
rect 2450 -585 2460 -115
rect 2480 -585 2490 -115
rect 2450 -595 2490 -585
rect 3700 -115 3740 -105
rect 3700 -585 3710 -115
rect 3730 -585 3740 -115
rect 3700 -595 3740 -585
<< end >>
