magic
tech sky130A
timestamp 1617765373
<< error_p >>
rect 6474 -112 6480 -109
rect 12974 -112 12980 -109
rect 6457 -115 6483 -112
rect 12957 -115 12983 -112
rect 6454 -118 6486 -115
rect 6454 -121 6463 -118
rect 6460 -582 6463 -121
rect 6477 -121 6486 -118
rect 12954 -118 12986 -115
rect 12954 -121 12963 -118
rect 6477 -582 6483 -121
rect 6460 -585 6483 -582
rect 12960 -582 12963 -121
rect 12977 -121 12986 -118
rect 12977 -582 12983 -121
rect 12960 -585 12983 -582
rect 6474 -588 6483 -585
rect 12974 -588 12983 -585
rect 6474 -591 6480 -588
rect 12974 -591 12980 -588
rect 4274 -927 4280 -924
rect 9724 -927 9730 -924
rect 4257 -930 4283 -927
rect 9707 -930 9733 -927
rect 4254 -933 4286 -930
rect 4254 -936 4263 -933
rect 4260 -1397 4263 -936
rect 4277 -936 4286 -933
rect 9704 -933 9736 -930
rect 9704 -936 9713 -933
rect 4277 -1397 4283 -936
rect 4260 -1400 4283 -1397
rect 9710 -1397 9713 -936
rect 9727 -936 9736 -933
rect 9727 -1397 9733 -936
rect 9710 -1400 9733 -1397
rect 4274 -1403 4283 -1400
rect 9724 -1403 9733 -1400
rect 4274 -1406 4280 -1403
rect 9724 -1406 9730 -1403
rect 6374 -1777 6380 -1774
rect 6424 -1777 6430 -1774
rect 6474 -1777 6480 -1774
rect 10774 -1777 10780 -1774
rect 10824 -1777 10830 -1774
rect 10874 -1777 10880 -1774
rect 6357 -1780 6383 -1777
rect 6407 -1780 6433 -1777
rect 6457 -1780 6483 -1777
rect 10757 -1780 10783 -1777
rect 10807 -1780 10833 -1777
rect 10857 -1780 10883 -1777
rect 6354 -1783 6386 -1780
rect 6354 -1786 6363 -1783
rect 6360 -2247 6363 -1786
rect 6377 -1786 6386 -1783
rect 6404 -1783 6436 -1780
rect 6404 -1786 6413 -1783
rect 6377 -2247 6383 -1786
rect 6360 -2250 6383 -2247
rect 6410 -2247 6413 -1786
rect 6427 -1786 6436 -1783
rect 6454 -1783 6486 -1780
rect 6454 -1786 6463 -1783
rect 6427 -2247 6433 -1786
rect 6410 -2250 6433 -2247
rect 6460 -2247 6463 -1786
rect 6477 -1786 6486 -1783
rect 10754 -1783 10786 -1780
rect 10754 -1786 10763 -1783
rect 6477 -2247 6483 -1786
rect 6460 -2250 6483 -2247
rect 10760 -2247 10763 -1786
rect 10777 -1786 10786 -1783
rect 10804 -1783 10836 -1780
rect 10804 -1786 10813 -1783
rect 10777 -2247 10783 -1786
rect 10760 -2250 10783 -2247
rect 10810 -2247 10813 -1786
rect 10827 -1786 10836 -1783
rect 10854 -1783 10886 -1780
rect 10854 -1786 10863 -1783
rect 10827 -2247 10833 -1786
rect 10810 -2250 10833 -2247
rect 10860 -2247 10863 -1786
rect 10877 -1786 10886 -1783
rect 10877 -2247 10883 -1786
rect 10860 -2250 10883 -2247
rect 6374 -2253 6383 -2250
rect 6424 -2253 6433 -2250
rect 6474 -2253 6483 -2250
rect 10774 -2253 10783 -2250
rect 10824 -2253 10833 -2250
rect 10874 -2253 10883 -2250
rect 6374 -2256 6380 -2253
rect 6424 -2256 6430 -2253
rect 6474 -2256 6480 -2253
rect 10774 -2256 10780 -2253
rect 10824 -2256 10830 -2253
rect 10874 -2256 10880 -2253
rect 6374 -2477 6380 -2474
rect 6424 -2477 6430 -2474
rect 6474 -2477 6480 -2474
rect 8574 -2477 8580 -2474
rect 8624 -2477 8630 -2474
rect 8674 -2477 8680 -2474
rect 10774 -2477 10780 -2474
rect 10824 -2477 10830 -2474
rect 10874 -2477 10880 -2474
rect 6357 -2480 6383 -2477
rect 6407 -2480 6433 -2477
rect 6457 -2480 6483 -2477
rect 8557 -2480 8583 -2477
rect 8607 -2480 8633 -2477
rect 8657 -2480 8683 -2477
rect 10757 -2480 10783 -2477
rect 10807 -2480 10833 -2477
rect 10857 -2480 10883 -2477
rect 6354 -2483 6386 -2480
rect 6354 -2486 6363 -2483
rect 6360 -2947 6363 -2486
rect 6377 -2486 6386 -2483
rect 6404 -2483 6436 -2480
rect 6404 -2486 6413 -2483
rect 6377 -2947 6383 -2486
rect 6360 -2950 6383 -2947
rect 6410 -2947 6413 -2486
rect 6427 -2486 6436 -2483
rect 6454 -2483 6486 -2480
rect 6454 -2486 6463 -2483
rect 6427 -2947 6433 -2486
rect 6410 -2950 6433 -2947
rect 6460 -2947 6463 -2486
rect 6477 -2486 6486 -2483
rect 8554 -2483 8586 -2480
rect 8554 -2486 8563 -2483
rect 6477 -2947 6483 -2486
rect 6460 -2950 6483 -2947
rect 8560 -2947 8563 -2486
rect 8577 -2486 8586 -2483
rect 8604 -2483 8636 -2480
rect 8604 -2486 8613 -2483
rect 8577 -2947 8583 -2486
rect 8560 -2950 8583 -2947
rect 8610 -2947 8613 -2486
rect 8627 -2486 8636 -2483
rect 8654 -2483 8686 -2480
rect 8654 -2486 8663 -2483
rect 8627 -2947 8633 -2486
rect 8610 -2950 8633 -2947
rect 8660 -2947 8663 -2486
rect 8677 -2486 8686 -2483
rect 10754 -2483 10786 -2480
rect 10754 -2486 10763 -2483
rect 8677 -2947 8683 -2486
rect 8660 -2950 8683 -2947
rect 10760 -2947 10763 -2486
rect 10777 -2486 10786 -2483
rect 10804 -2483 10836 -2480
rect 10804 -2486 10813 -2483
rect 10777 -2947 10783 -2486
rect 10760 -2950 10783 -2947
rect 10810 -2947 10813 -2486
rect 10827 -2486 10836 -2483
rect 10854 -2483 10886 -2480
rect 10854 -2486 10863 -2483
rect 10827 -2947 10833 -2486
rect 10810 -2950 10833 -2947
rect 10860 -2947 10863 -2486
rect 10877 -2486 10886 -2483
rect 10877 -2947 10883 -2486
rect 10860 -2950 10883 -2947
rect 6374 -2953 6383 -2950
rect 6424 -2953 6433 -2950
rect 6474 -2953 6483 -2950
rect 8574 -2953 8583 -2950
rect 8624 -2953 8633 -2950
rect 8674 -2953 8683 -2950
rect 10774 -2953 10783 -2950
rect 10824 -2953 10833 -2950
rect 10874 -2953 10883 -2950
rect 6374 -2956 6380 -2953
rect 6424 -2956 6430 -2953
rect 6474 -2956 6480 -2953
rect 8574 -2956 8580 -2953
rect 8624 -2956 8630 -2953
rect 8674 -2956 8680 -2953
rect 10774 -2956 10780 -2953
rect 10824 -2956 10830 -2953
rect 10874 -2956 10880 -2953
<< nmos >>
rect -5 -600 995 -100
rect 1045 -600 2045 -100
rect 2195 -600 3195 -100
rect 3245 -600 4245 -100
rect 4295 -600 5295 -100
rect 5445 -600 6445 -100
rect 6495 -600 7495 -100
rect 7545 -600 8545 -100
rect 8695 -600 9695 -100
rect 9745 -600 10745 -100
rect 10895 -600 11895 -100
rect 11945 -600 12945 -100
rect 12995 -600 13995 -100
rect 14145 -600 15145 -100
rect -5 -1415 995 -915
rect 1045 -1415 2045 -915
rect 2195 -1415 3195 -915
rect 3245 -1415 4245 -915
rect 4295 -1415 5295 -915
rect 5445 -1415 6445 -915
rect 6495 -1415 7495 -915
rect 7545 -1415 8545 -915
rect 8695 -1415 9695 -915
rect 9745 -1415 10745 -915
rect 10795 -1415 11795 -915
rect 11945 -1415 12945 -915
rect 12995 -1415 13995 -915
rect 14145 -1415 15145 -915
rect 15195 -1415 16195 -915
rect 16345 -1415 17345 -915
rect 17395 -1415 18395 -915
rect 3245 -2265 4245 -1765
rect 4295 -2265 5295 -1765
rect 5345 -2265 6345 -1765
rect 6495 -2265 7495 -1765
rect 7545 -2265 8545 -1765
rect 8695 -2265 9695 -1765
rect 9745 -2265 10745 -1765
rect 10895 -2265 11895 -1765
rect 11945 -2265 12945 -1765
rect 12995 -2265 13995 -1765
rect 3245 -2965 4245 -2465
rect 4295 -2965 5295 -2465
rect 5345 -2965 6345 -2465
rect 6495 -2965 7495 -2465
rect 7545 -2965 8545 -2465
rect 8695 -2965 9695 -2465
rect 9745 -2965 10745 -2465
rect 10895 -2965 11895 -2465
rect 11945 -2965 12945 -2465
rect 12995 -2965 13995 -2465
<< ndiff >>
rect -55 -115 -5 -100
rect -55 -585 -40 -115
rect -20 -585 -5 -115
rect -55 -600 -5 -585
rect 995 -115 1045 -100
rect 995 -585 1010 -115
rect 1030 -585 1045 -115
rect 995 -600 1045 -585
rect 2045 -115 2095 -100
rect 2145 -115 2195 -100
rect 2045 -585 2060 -115
rect 2080 -585 2095 -115
rect 2145 -585 2160 -115
rect 2180 -585 2195 -115
rect 2045 -600 2095 -585
rect 2145 -600 2195 -585
rect 3195 -115 3245 -100
rect 3195 -585 3210 -115
rect 3230 -585 3245 -115
rect 3195 -600 3245 -585
rect 4245 -115 4295 -100
rect 4245 -585 4260 -115
rect 4280 -585 4295 -115
rect 4245 -600 4295 -585
rect 5295 -115 5345 -100
rect 5395 -115 5445 -100
rect 5295 -585 5310 -115
rect 5330 -585 5345 -115
rect 5395 -585 5410 -115
rect 5430 -585 5445 -115
rect 5295 -600 5345 -585
rect 5395 -600 5445 -585
rect 6445 -115 6495 -100
rect 6445 -585 6460 -115
rect 6480 -585 6495 -115
rect 6445 -600 6495 -585
rect 7495 -115 7545 -100
rect 7495 -585 7510 -115
rect 7530 -585 7545 -115
rect 7495 -600 7545 -585
rect 8545 -115 8595 -100
rect 8645 -115 8695 -100
rect 8545 -585 8560 -115
rect 8580 -585 8595 -115
rect 8645 -585 8660 -115
rect 8680 -585 8695 -115
rect 8545 -600 8595 -585
rect 8645 -600 8695 -585
rect 9695 -115 9745 -100
rect 9695 -585 9710 -115
rect 9730 -585 9745 -115
rect 9695 -600 9745 -585
rect 10745 -110 10795 -100
rect 10845 -110 10895 -100
rect 10745 -585 10760 -110
rect 10780 -585 10795 -110
rect 10845 -585 10860 -110
rect 10880 -585 10895 -110
rect 10745 -600 10795 -585
rect 10845 -600 10895 -585
rect 11895 -115 11945 -100
rect 11895 -585 11910 -115
rect 11930 -585 11945 -115
rect 11895 -600 11945 -585
rect 12945 -115 12995 -100
rect 12945 -585 12960 -115
rect 12980 -585 12995 -115
rect 12945 -600 12995 -585
rect 13995 -115 14045 -100
rect 14095 -115 14145 -100
rect 13995 -585 14010 -115
rect 14030 -585 14045 -115
rect 14095 -585 14110 -115
rect 14130 -585 14145 -115
rect 13995 -600 14045 -585
rect 14095 -600 14145 -585
rect 15145 -115 15195 -100
rect 15145 -585 15160 -115
rect 15180 -585 15195 -115
rect 15145 -600 15195 -585
rect -55 -930 -5 -915
rect -55 -1400 -40 -930
rect -20 -1400 -5 -930
rect -55 -1415 -5 -1400
rect 995 -930 1045 -915
rect 995 -1400 1010 -930
rect 1030 -1400 1045 -930
rect 995 -1415 1045 -1400
rect 2045 -930 2095 -915
rect 2145 -930 2195 -915
rect 2045 -1400 2060 -930
rect 2080 -1400 2095 -930
rect 2145 -1400 2160 -930
rect 2180 -1400 2195 -930
rect 2045 -1415 2095 -1400
rect 2145 -1415 2195 -1400
rect 3195 -930 3245 -915
rect 3195 -1400 3210 -930
rect 3230 -1400 3245 -930
rect 3195 -1415 3245 -1400
rect 4245 -930 4295 -915
rect 4245 -1400 4260 -930
rect 4280 -1400 4295 -930
rect 4245 -1415 4295 -1400
rect 5295 -930 5345 -915
rect 5395 -930 5445 -915
rect 5295 -1400 5310 -930
rect 5330 -1400 5345 -930
rect 5395 -1400 5410 -930
rect 5430 -1400 5445 -930
rect 5295 -1415 5345 -1400
rect 5395 -1415 5445 -1400
rect 6445 -930 6495 -915
rect 6445 -1400 6460 -930
rect 6480 -1400 6495 -930
rect 6445 -1415 6495 -1400
rect 7495 -930 7545 -915
rect 7495 -1400 7510 -930
rect 7530 -1400 7545 -930
rect 7495 -1415 7545 -1400
rect 8545 -930 8595 -915
rect 8645 -930 8695 -915
rect 8545 -1400 8560 -930
rect 8580 -1400 8595 -930
rect 8645 -1400 8660 -930
rect 8680 -1400 8695 -930
rect 8545 -1415 8595 -1400
rect 8645 -1415 8695 -1400
rect 9695 -930 9745 -915
rect 9695 -1400 9710 -930
rect 9730 -1400 9745 -930
rect 9695 -1415 9745 -1400
rect 10745 -930 10795 -915
rect 10745 -1400 10760 -930
rect 10780 -1400 10795 -930
rect 10745 -1415 10795 -1400
rect 11795 -930 11845 -915
rect 11895 -930 11945 -915
rect 11795 -1400 11810 -930
rect 11830 -1400 11845 -930
rect 11895 -1400 11910 -930
rect 11930 -1400 11945 -930
rect 11795 -1415 11845 -1400
rect 11895 -1415 11945 -1400
rect 12945 -930 12995 -915
rect 12945 -1400 12960 -930
rect 12980 -1400 12995 -930
rect 12945 -1415 12995 -1400
rect 13995 -930 14045 -915
rect 14095 -930 14145 -915
rect 13995 -1400 14010 -930
rect 14030 -1400 14045 -930
rect 14095 -1400 14110 -930
rect 14130 -1400 14145 -930
rect 13995 -1415 14045 -1400
rect 14095 -1415 14145 -1400
rect 15145 -930 15195 -915
rect 15145 -1400 15160 -930
rect 15180 -1400 15195 -930
rect 15145 -1415 15195 -1400
rect 16195 -930 16245 -915
rect 16295 -930 16345 -915
rect 16195 -1400 16210 -930
rect 16230 -1400 16245 -930
rect 16295 -1400 16310 -930
rect 16330 -1400 16345 -930
rect 16195 -1415 16245 -1400
rect 16295 -1415 16345 -1400
rect 17345 -930 17395 -915
rect 17345 -1400 17360 -930
rect 17380 -1400 17395 -930
rect 17345 -1415 17395 -1400
rect 18395 -930 18445 -915
rect 18395 -1400 18410 -930
rect 18430 -1400 18445 -930
rect 18395 -1415 18445 -1400
rect 3195 -1780 3245 -1765
rect 3195 -2250 3210 -1780
rect 3230 -2250 3245 -1780
rect 3195 -2265 3245 -2250
rect 4245 -1780 4295 -1765
rect 4245 -2250 4260 -1780
rect 4280 -2250 4295 -1780
rect 4245 -2265 4295 -2250
rect 5295 -1780 5345 -1765
rect 5295 -2250 5310 -1780
rect 5330 -2250 5345 -1780
rect 5295 -2265 5345 -2250
rect 6345 -1780 6395 -1765
rect 6445 -1780 6495 -1765
rect 6345 -2250 6360 -1780
rect 6380 -2250 6395 -1780
rect 6445 -2250 6460 -1780
rect 6480 -2250 6495 -1780
rect 6345 -2265 6395 -2250
rect 6445 -2265 6495 -2250
rect 7495 -1780 7545 -1765
rect 7495 -2250 7510 -1780
rect 7530 -2250 7545 -1780
rect 7495 -2265 7545 -2250
rect 8545 -1780 8595 -1765
rect 8645 -1780 8695 -1765
rect 8545 -2250 8560 -1780
rect 8580 -2250 8595 -1780
rect 8645 -2250 8660 -1780
rect 8680 -2250 8695 -1780
rect 8545 -2265 8595 -2250
rect 8645 -2265 8695 -2250
rect 9695 -1780 9745 -1765
rect 9695 -2250 9710 -1780
rect 9730 -2250 9745 -1780
rect 9695 -2265 9745 -2250
rect 10745 -1780 10795 -1765
rect 10845 -1780 10895 -1765
rect 10745 -2250 10760 -1780
rect 10780 -2250 10795 -1780
rect 10845 -2250 10860 -1780
rect 10880 -2250 10895 -1780
rect 10745 -2265 10795 -2250
rect 10845 -2265 10895 -2250
rect 11895 -1780 11945 -1765
rect 11895 -2250 11910 -1780
rect 11930 -2250 11945 -1780
rect 11895 -2265 11945 -2250
rect 12945 -1780 12995 -1765
rect 12945 -2250 12960 -1780
rect 12980 -2250 12995 -1780
rect 12945 -2265 12995 -2250
rect 13995 -1780 14045 -1765
rect 13995 -2250 14010 -1780
rect 14030 -2250 14045 -1780
rect 13995 -2265 14045 -2250
rect 3195 -2480 3245 -2465
rect 3195 -2950 3210 -2480
rect 3230 -2950 3245 -2480
rect 3195 -2965 3245 -2950
rect 4245 -2480 4295 -2465
rect 4245 -2950 4260 -2480
rect 4280 -2950 4295 -2480
rect 4245 -2965 4295 -2950
rect 5295 -2480 5345 -2465
rect 5295 -2950 5310 -2480
rect 5330 -2950 5345 -2480
rect 5295 -2965 5345 -2950
rect 6345 -2480 6395 -2465
rect 6445 -2480 6495 -2465
rect 6345 -2950 6360 -2480
rect 6380 -2950 6395 -2480
rect 6445 -2950 6460 -2480
rect 6480 -2950 6495 -2480
rect 6345 -2965 6395 -2950
rect 6445 -2965 6495 -2950
rect 7495 -2480 7545 -2465
rect 7495 -2950 7510 -2480
rect 7530 -2950 7545 -2480
rect 7495 -2965 7545 -2950
rect 8545 -2480 8595 -2465
rect 8645 -2480 8695 -2465
rect 8545 -2950 8560 -2480
rect 8580 -2950 8595 -2480
rect 8645 -2950 8660 -2480
rect 8680 -2950 8695 -2480
rect 8545 -2965 8595 -2950
rect 8645 -2965 8695 -2950
rect 9695 -2480 9745 -2465
rect 9695 -2950 9710 -2480
rect 9730 -2950 9745 -2480
rect 9695 -2965 9745 -2950
rect 10745 -2480 10795 -2465
rect 10845 -2480 10895 -2465
rect 10745 -2950 10760 -2480
rect 10780 -2950 10795 -2480
rect 10845 -2950 10860 -2480
rect 10880 -2950 10895 -2480
rect 10745 -2965 10795 -2950
rect 10845 -2965 10895 -2950
rect 11895 -2480 11945 -2465
rect 11895 -2950 11910 -2480
rect 11930 -2950 11945 -2480
rect 11895 -2965 11945 -2950
rect 12945 -2480 12995 -2465
rect 12945 -2950 12960 -2480
rect 12980 -2950 12995 -2480
rect 12945 -2965 12995 -2950
rect 13995 -2480 14045 -2465
rect 13995 -2950 14010 -2480
rect 14030 -2950 14045 -2480
rect 13995 -2965 14045 -2950
<< ndiffc >>
rect -40 -585 -20 -115
rect 1010 -585 1030 -115
rect 2060 -585 2080 -115
rect 2160 -585 2180 -115
rect 3210 -585 3230 -115
rect 4260 -585 4280 -115
rect 5310 -585 5330 -115
rect 5410 -585 5430 -115
rect 6460 -585 6480 -115
rect 7510 -585 7530 -115
rect 8560 -585 8580 -115
rect 8660 -585 8680 -115
rect 9710 -585 9730 -115
rect 10760 -585 10780 -110
rect 10860 -585 10880 -110
rect 11910 -585 11930 -115
rect 12960 -585 12980 -115
rect 14010 -585 14030 -115
rect 14110 -585 14130 -115
rect 15160 -585 15180 -115
rect -40 -1400 -20 -930
rect 1010 -1400 1030 -930
rect 2060 -1400 2080 -930
rect 2160 -1400 2180 -930
rect 3210 -1400 3230 -930
rect 4260 -1400 4280 -930
rect 5310 -1400 5330 -930
rect 5410 -1400 5430 -930
rect 6460 -1400 6480 -930
rect 7510 -1400 7530 -930
rect 8560 -1400 8580 -930
rect 8660 -1400 8680 -930
rect 9710 -1400 9730 -930
rect 10760 -1400 10780 -930
rect 11810 -1400 11830 -930
rect 11910 -1400 11930 -930
rect 12960 -1400 12980 -930
rect 14010 -1400 14030 -930
rect 14110 -1400 14130 -930
rect 15160 -1400 15180 -930
rect 16210 -1400 16230 -930
rect 16310 -1400 16330 -930
rect 17360 -1400 17380 -930
rect 18410 -1400 18430 -930
rect 3210 -2250 3230 -1780
rect 4260 -2250 4280 -1780
rect 5310 -2250 5330 -1780
rect 6360 -2250 6380 -1780
rect 6460 -2250 6480 -1780
rect 7510 -2250 7530 -1780
rect 8560 -2250 8580 -1780
rect 8660 -2250 8680 -1780
rect 9710 -2250 9730 -1780
rect 10760 -2250 10780 -1780
rect 10860 -2250 10880 -1780
rect 11910 -2250 11930 -1780
rect 12960 -2250 12980 -1780
rect 14010 -2250 14030 -1780
rect 3210 -2950 3230 -2480
rect 4260 -2950 4280 -2480
rect 5310 -2950 5330 -2480
rect 6360 -2950 6380 -2480
rect 6460 -2950 6480 -2480
rect 7510 -2950 7530 -2480
rect 8560 -2950 8580 -2480
rect 8660 -2950 8680 -2480
rect 9710 -2950 9730 -2480
rect 10760 -2950 10780 -2480
rect 10860 -2950 10880 -2480
rect 11910 -2950 11930 -2480
rect 12960 -2950 12980 -2480
rect 14010 -2950 14030 -2480
<< psubdiff >>
rect -105 -115 -55 -100
rect -105 -585 -90 -115
rect -70 -585 -55 -115
rect -105 -600 -55 -585
rect 2095 -115 2145 -100
rect 2095 -585 2110 -115
rect 2130 -585 2145 -115
rect 2095 -600 2145 -585
rect 5345 -115 5395 -100
rect 5345 -585 5360 -115
rect 5380 -585 5395 -115
rect 5345 -600 5395 -585
rect 8595 -115 8645 -100
rect 8595 -585 8610 -115
rect 8630 -585 8645 -115
rect 8595 -600 8645 -585
rect 10795 -110 10845 -100
rect 10795 -585 10810 -110
rect 10830 -585 10845 -110
rect 10795 -600 10845 -585
rect 14045 -115 14095 -100
rect 14045 -585 14060 -115
rect 14080 -585 14095 -115
rect 14045 -600 14095 -585
rect -105 -930 -55 -915
rect -105 -1400 -90 -930
rect -70 -1400 -55 -930
rect -105 -1415 -55 -1400
rect 2095 -930 2145 -915
rect 2095 -1400 2110 -930
rect 2130 -1400 2145 -930
rect 2095 -1415 2145 -1400
rect 5345 -930 5395 -915
rect 5345 -1400 5360 -930
rect 5380 -1400 5395 -930
rect 5345 -1415 5395 -1400
rect 8595 -930 8645 -915
rect 8595 -1400 8610 -930
rect 8630 -1400 8645 -930
rect 8595 -1415 8645 -1400
rect 11845 -930 11895 -915
rect 11845 -1400 11860 -930
rect 11880 -1400 11895 -930
rect 11845 -1415 11895 -1400
rect 14045 -930 14095 -915
rect 14045 -1400 14060 -930
rect 14080 -1400 14095 -930
rect 14045 -1415 14095 -1400
rect 16245 -930 16295 -915
rect 16245 -1400 16260 -930
rect 16280 -1400 16295 -930
rect 16245 -1415 16295 -1400
rect 18445 -930 18495 -915
rect 18445 -1400 18460 -930
rect 18480 -1400 18495 -930
rect 18445 -1415 18495 -1400
rect 3145 -1780 3195 -1765
rect 3145 -2250 3160 -1780
rect 3180 -2250 3195 -1780
rect 3145 -2265 3195 -2250
rect 6395 -1780 6445 -1765
rect 6395 -2250 6410 -1780
rect 6430 -2250 6445 -1780
rect 6395 -2265 6445 -2250
rect 8595 -1780 8645 -1765
rect 8595 -2250 8610 -1780
rect 8630 -2250 8645 -1780
rect 8595 -2265 8645 -2250
rect 10795 -1780 10845 -1765
rect 10795 -2250 10810 -1780
rect 10830 -2250 10845 -1780
rect 10795 -2265 10845 -2250
rect 14045 -1780 14095 -1765
rect 14045 -2250 14060 -1780
rect 14080 -2250 14095 -1780
rect 14045 -2265 14095 -2250
rect 3145 -2480 3195 -2465
rect 3145 -2950 3160 -2480
rect 3180 -2950 3195 -2480
rect 3145 -2965 3195 -2950
rect 6395 -2480 6445 -2465
rect 6395 -2950 6410 -2480
rect 6430 -2950 6445 -2480
rect 6395 -2965 6445 -2950
rect 8595 -2480 8645 -2465
rect 8595 -2950 8610 -2480
rect 8630 -2950 8645 -2480
rect 8595 -2965 8645 -2950
rect 10795 -2480 10845 -2465
rect 10795 -2950 10810 -2480
rect 10830 -2950 10845 -2480
rect 10795 -2965 10845 -2950
rect 14045 -2480 14095 -2465
rect 14045 -2950 14060 -2480
rect 14080 -2950 14095 -2480
rect 14045 -2965 14095 -2950
<< psubdiffcont >>
rect -90 -585 -70 -115
rect 2110 -585 2130 -115
rect 5360 -585 5380 -115
rect 8610 -585 8630 -115
rect 10810 -585 10830 -110
rect 14060 -585 14080 -115
rect -90 -1400 -70 -930
rect 2110 -1400 2130 -930
rect 5360 -1400 5380 -930
rect 8610 -1400 8630 -930
rect 11860 -1400 11880 -930
rect 14060 -1400 14080 -930
rect 16260 -1400 16280 -930
rect 18460 -1400 18480 -930
rect 3160 -2250 3180 -1780
rect 6410 -2250 6430 -1780
rect 8610 -2250 8630 -1780
rect 10810 -2250 10830 -1780
rect 14060 -2250 14080 -1780
rect 3160 -2950 3180 -2480
rect 6410 -2950 6430 -2480
rect 8610 -2950 8630 -2480
rect 10810 -2950 10830 -2480
rect 14060 -2950 14080 -2480
<< poly >>
rect 1045 -45 13995 -30
rect -50 -55 -10 -45
rect -50 -75 -40 -55
rect -20 -70 -10 -55
rect -20 -75 995 -70
rect -50 -85 995 -75
rect -5 -100 995 -85
rect 1045 -100 2045 -45
rect 2195 -100 3195 -45
rect 3245 -100 4245 -45
rect 4295 -100 5295 -45
rect 5445 -100 6445 -45
rect 6495 -100 7495 -45
rect 7545 -100 8545 -70
rect 8695 -100 9695 -70
rect 9745 -100 10745 -45
rect 10895 -100 11895 -45
rect 11945 -100 12945 -45
rect 12995 -100 13995 -45
rect 15150 -55 15190 -45
rect 15150 -70 15160 -55
rect 14145 -75 15160 -70
rect 15180 -75 15190 -55
rect 14145 -85 15190 -75
rect 14145 -100 15145 -85
rect -5 -615 995 -600
rect 1045 -615 2045 -600
rect 2195 -615 3195 -600
rect 3245 -615 4245 -600
rect 4295 -615 5295 -600
rect 5445 -615 6445 -600
rect 6495 -615 7495 -600
rect 7545 -615 8545 -600
rect 8695 -615 9695 -600
rect 9745 -615 10745 -600
rect 10895 -615 11895 -600
rect 11945 -615 12945 -600
rect 12995 -615 13995 -600
rect 14145 -615 15145 -600
rect 1045 -745 1090 -615
rect 7545 -625 9695 -615
rect 7545 -630 8610 -625
rect 2005 -650 2045 -640
rect 2195 -650 2235 -640
rect 2005 -670 2015 -650
rect 2035 -670 2205 -650
rect 2225 -670 2235 -650
rect 2005 -680 2045 -670
rect 2195 -680 2235 -670
rect 4190 -650 4230 -640
rect 4310 -650 4350 -640
rect 4190 -670 4200 -650
rect 4220 -670 4320 -650
rect 4340 -670 4350 -650
rect 8600 -645 8610 -630
rect 8630 -630 9695 -625
rect 8630 -645 8640 -630
rect 8600 -655 8640 -645
rect 10685 -650 10725 -640
rect 10915 -650 10955 -640
rect 4190 -680 4230 -670
rect 4310 -680 4350 -670
rect 10685 -670 10695 -650
rect 10715 -670 10925 -650
rect 10945 -670 10955 -650
rect 10685 -680 10725 -670
rect 10915 -680 10955 -670
rect 8480 -710 8520 -700
rect 8720 -710 8760 -700
rect 8480 -730 8490 -710
rect 8510 -730 8730 -710
rect 8750 -730 8760 -710
rect 8480 -740 8520 -730
rect 8720 -740 8760 -730
rect 1045 -770 1055 -745
rect 1080 -770 1090 -745
rect 1045 -860 1090 -770
rect -50 -870 -10 -860
rect -50 -890 -40 -870
rect -20 -885 -10 -870
rect 1045 -875 17345 -860
rect -20 -890 995 -885
rect -50 -900 995 -890
rect -5 -915 995 -900
rect 1045 -915 2045 -875
rect 2195 -915 3195 -875
rect 3245 -915 4245 -875
rect 4295 -915 5295 -875
rect 5445 -915 6445 -875
rect 6495 -915 7495 -875
rect 7545 -915 8545 -900
rect 8695 -915 9695 -900
rect 9745 -915 10745 -875
rect 10795 -915 11795 -875
rect 11945 -915 12945 -875
rect 12995 -915 13995 -900
rect 14145 -915 15145 -900
rect 15195 -915 16195 -875
rect 16345 -915 17345 -875
rect 18455 -870 18495 -860
rect 18455 -885 18465 -870
rect 17395 -890 18465 -885
rect 18485 -890 18495 -870
rect 17395 -900 18495 -890
rect 17395 -915 18395 -900
rect -5 -1430 995 -1415
rect 1045 -1430 2045 -1415
rect 2195 -1430 3195 -1415
rect 3245 -1430 4245 -1415
rect 4295 -1430 5295 -1415
rect 5445 -1430 6445 -1415
rect 6495 -1430 7495 -1415
rect 7545 -1430 8545 -1415
rect 8695 -1430 9695 -1415
rect 9745 -1430 10745 -1415
rect 10795 -1430 11795 -1415
rect 11945 -1430 12945 -1415
rect 12995 -1430 13995 -1415
rect 14145 -1430 15145 -1415
rect 15195 -1430 16195 -1415
rect 16345 -1430 17345 -1415
rect 17395 -1430 18395 -1415
rect 1045 -1505 1090 -1430
rect 7545 -1440 9695 -1430
rect 7545 -1445 8610 -1440
rect 2005 -1465 2045 -1455
rect 2195 -1465 2235 -1455
rect 2005 -1485 2015 -1465
rect 2035 -1485 2205 -1465
rect 2225 -1485 2235 -1465
rect 8600 -1460 8610 -1445
rect 8630 -1445 9695 -1440
rect 12995 -1440 15145 -1430
rect 12995 -1445 14060 -1440
rect 8630 -1460 8640 -1445
rect 8600 -1470 8640 -1460
rect 14050 -1460 14060 -1445
rect 14080 -1445 15145 -1440
rect 14080 -1460 14090 -1445
rect 14050 -1470 14090 -1460
rect 2005 -1495 2045 -1485
rect 2195 -1495 2235 -1485
rect 12875 -1500 12915 -1490
rect 13025 -1500 13065 -1490
rect 6355 -1525 6395 -1515
rect 6545 -1525 6585 -1515
rect 6355 -1545 6365 -1525
rect 6385 -1545 6555 -1525
rect 6575 -1545 6585 -1525
rect 12875 -1520 12885 -1500
rect 12905 -1520 13035 -1500
rect 13055 -1520 13065 -1500
rect 12875 -1530 12915 -1520
rect 13025 -1530 13065 -1520
rect 6355 -1555 6395 -1545
rect 6545 -1555 6585 -1545
rect 8535 -1585 8575 -1575
rect 8665 -1585 8705 -1575
rect 2005 -1610 2045 -1600
rect 2195 -1610 2235 -1600
rect 2005 -1630 2015 -1610
rect 2035 -1630 2205 -1610
rect 2225 -1630 2235 -1610
rect 8535 -1605 8545 -1585
rect 8565 -1605 8675 -1585
rect 8695 -1605 8705 -1585
rect 8535 -1615 8575 -1605
rect 8665 -1615 8705 -1605
rect 2005 -1640 2045 -1630
rect 2195 -1640 2235 -1630
rect 2005 -1675 2045 -1665
rect 2195 -1675 2235 -1665
rect 2005 -1695 2015 -1675
rect 2035 -1695 2205 -1675
rect 2225 -1695 2235 -1675
rect 2005 -1705 2045 -1695
rect 2195 -1705 2235 -1695
rect 3245 -1765 4245 -1750
rect 4295 -1765 5295 -1750
rect 5345 -1765 6345 -1750
rect 6495 -1765 7495 -1750
rect 7545 -1765 8545 -1750
rect 8695 -1765 9695 -1750
rect 9745 -1765 10745 -1750
rect 10895 -1765 11895 -1750
rect 11945 -1765 12945 -1750
rect 12995 -1765 13995 -1750
rect 3245 -2280 4245 -2265
rect 4295 -2280 5295 -2265
rect 5345 -2280 6345 -2265
rect 6495 -2280 7495 -2265
rect 7545 -2280 8545 -2265
rect 8695 -2280 9695 -2265
rect 9745 -2280 10745 -2265
rect 10895 -2280 11895 -2265
rect 11945 -2280 12945 -2265
rect 12995 -2280 13995 -2265
rect 7545 -2290 9695 -2280
rect 7545 -2295 8610 -2290
rect 8600 -2310 8610 -2295
rect 8630 -2295 9695 -2290
rect 8630 -2310 8640 -2295
rect 8600 -2320 8640 -2310
rect 3245 -2465 4245 -2450
rect 4295 -2465 5295 -2450
rect 5345 -2465 6345 -2450
rect 6495 -2465 7495 -2450
rect 7545 -2465 8545 -2450
rect 8695 -2465 9695 -2450
rect 9745 -2465 10745 -2450
rect 10895 -2465 11895 -2450
rect 11945 -2465 12945 -2450
rect 12995 -2465 13995 -2450
rect 3245 -2980 4245 -2965
rect 4295 -2980 5295 -2965
rect 5345 -2980 6345 -2965
rect 6495 -2980 7495 -2965
rect 7545 -2980 8545 -2965
rect 8695 -2980 9695 -2965
rect 9745 -2980 10745 -2965
rect 10895 -2980 11895 -2965
rect 11945 -2980 12945 -2965
rect 12995 -2980 13995 -2965
rect 7545 -2990 9695 -2980
rect 7545 -2995 8610 -2990
rect 8600 -3010 8610 -2995
rect 8630 -2995 9695 -2990
rect 8630 -3010 8640 -2995
rect 8600 -3020 8640 -3010
<< polycont >>
rect -40 -75 -20 -55
rect 15160 -75 15180 -55
rect 2015 -670 2035 -650
rect 2205 -670 2225 -650
rect 4200 -670 4220 -650
rect 4320 -670 4340 -650
rect 8610 -645 8630 -625
rect 10695 -670 10715 -650
rect 10925 -670 10945 -650
rect 8490 -730 8510 -710
rect 8730 -730 8750 -710
rect 1055 -770 1080 -745
rect -40 -890 -20 -870
rect 18465 -890 18485 -870
rect 2015 -1485 2035 -1465
rect 2205 -1485 2225 -1465
rect 8610 -1460 8630 -1440
rect 14060 -1460 14080 -1440
rect 6365 -1545 6385 -1525
rect 6555 -1545 6575 -1525
rect 12885 -1520 12905 -1500
rect 13035 -1520 13055 -1500
rect 2015 -1630 2035 -1610
rect 2205 -1630 2225 -1610
rect 8545 -1605 8565 -1585
rect 8675 -1605 8695 -1585
rect 2015 -1695 2035 -1675
rect 2205 -1695 2225 -1675
rect 8610 -2310 8630 -2290
rect 8610 -3010 8630 -2990
<< locali >>
rect -50 -55 -10 -45
rect -50 -75 -40 -55
rect -20 -75 -10 -55
rect -50 -105 -10 -75
rect 15150 -55 15190 -45
rect 15150 -75 15160 -55
rect 15180 -75 15190 -55
rect 15150 -105 15190 -75
rect -100 -115 -10 -105
rect -100 -585 -90 -115
rect -70 -585 -40 -115
rect -20 -585 -10 -115
rect -100 -595 -10 -585
rect 1000 -115 1040 -105
rect 1000 -585 1010 -115
rect 1030 -585 1040 -115
rect 1000 -640 1040 -585
rect 2050 -115 2190 -105
rect 2050 -585 2060 -115
rect 2080 -585 2110 -115
rect 2130 -585 2160 -115
rect 2180 -585 2190 -115
rect 2050 -595 2190 -585
rect 3200 -115 3240 -105
rect 3200 -585 3210 -115
rect 3230 -585 3240 -115
rect 1000 -650 2045 -640
rect 1000 -670 2015 -650
rect 2035 -670 2045 -650
rect 1000 -680 2045 -670
rect 2100 -700 2140 -595
rect 3200 -640 3240 -585
rect 4250 -115 4290 -105
rect 4250 -585 4260 -115
rect 4280 -585 4290 -115
rect 2195 -650 4230 -640
rect 2195 -670 2205 -650
rect 2225 -670 4200 -650
rect 4220 -670 4230 -650
rect 2195 -680 4230 -670
rect 4250 -700 4290 -585
rect 5300 -115 5440 -105
rect 5300 -585 5310 -115
rect 5330 -585 5360 -115
rect 5380 -585 5410 -115
rect 5430 -585 5440 -115
rect 5300 -595 5440 -585
rect 6450 -115 6490 -105
rect 6450 -585 6460 -115
rect 6480 -585 6490 -115
rect 6450 -595 6490 -585
rect 7500 -115 7540 -105
rect 7500 -585 7510 -115
rect 7530 -585 7540 -115
rect 5350 -640 5390 -595
rect 4310 -650 5390 -640
rect 4310 -670 4320 -650
rect 4340 -670 5390 -650
rect 4310 -680 5390 -670
rect 7500 -700 7540 -585
rect 8550 -115 8690 -105
rect 8550 -585 8560 -115
rect 8580 -585 8610 -115
rect 8630 -585 8660 -115
rect 8680 -585 8690 -115
rect 8550 -595 8690 -585
rect 9700 -115 9740 -105
rect 9700 -585 9710 -115
rect 9730 -585 9740 -115
rect 8605 -615 8635 -595
rect 8600 -625 8640 -615
rect 8600 -645 8610 -625
rect 8630 -645 8640 -625
rect 8600 -655 8640 -645
rect 9700 -640 9740 -585
rect 10750 -110 10890 -105
rect 10750 -585 10760 -110
rect 10780 -585 10810 -110
rect 10830 -585 10860 -110
rect 10880 -585 10890 -110
rect 10750 -595 10890 -585
rect 11900 -115 11940 -105
rect 11900 -585 11910 -115
rect 11930 -585 11940 -115
rect 9700 -650 10725 -640
rect -380 -745 1090 -735
rect -380 -770 1055 -745
rect 1080 -770 1090 -745
rect -380 -780 1090 -770
rect 1170 -740 3240 -700
rect 4250 -710 8520 -700
rect 4250 -730 8490 -710
rect 8510 -730 8520 -710
rect 4250 -740 8520 -730
rect 1170 -800 1210 -740
rect -180 -840 1210 -800
rect -180 -1665 -140 -840
rect -50 -870 -10 -860
rect -50 -890 -40 -870
rect -20 -890 -10 -870
rect -50 -920 -10 -890
rect -100 -930 -10 -920
rect -100 -1400 -90 -930
rect -70 -1400 -40 -930
rect -20 -1400 -10 -930
rect -100 -1410 -10 -1400
rect 1000 -930 1040 -920
rect 1000 -1400 1010 -930
rect 1030 -1400 1040 -930
rect 1000 -1455 1040 -1400
rect 2050 -930 2190 -920
rect 2050 -1400 2060 -930
rect 2080 -1400 2110 -930
rect 2130 -1400 2160 -930
rect 2180 -1400 2190 -930
rect 2050 -1410 2190 -1400
rect 3200 -930 3240 -740
rect 8605 -920 8635 -655
rect 9700 -670 10695 -650
rect 10715 -670 10725 -650
rect 9700 -680 10725 -670
rect 10800 -700 10840 -595
rect 11900 -640 11940 -585
rect 12950 -115 12990 -105
rect 12950 -585 12960 -115
rect 12980 -585 12990 -115
rect 12950 -595 12990 -585
rect 14000 -115 14140 -105
rect 14000 -585 14010 -115
rect 14030 -585 14060 -115
rect 14080 -585 14110 -115
rect 14130 -585 14140 -115
rect 14000 -595 14140 -585
rect 15145 -115 15190 -105
rect 15145 -585 15160 -115
rect 15180 -585 15190 -115
rect 15145 -595 15190 -585
rect 14050 -640 14090 -595
rect 10915 -650 18590 -640
rect 10915 -670 10925 -650
rect 10945 -670 18590 -650
rect 10915 -680 18590 -670
rect 8720 -710 10840 -700
rect 8720 -730 8730 -710
rect 8750 -730 10840 -710
rect 8720 -740 10840 -730
rect 16250 -850 16340 -810
rect 16250 -920 16290 -850
rect 18455 -870 18495 -860
rect 18455 -890 18465 -870
rect 18485 -890 18495 -870
rect 18455 -900 18495 -890
rect 18460 -920 18490 -900
rect 3200 -1400 3210 -930
rect 3230 -1400 3240 -930
rect 1000 -1465 2045 -1455
rect 1000 -1485 2015 -1465
rect 2035 -1485 2045 -1465
rect 1000 -1495 2045 -1485
rect 1000 -1600 1040 -1495
rect 2100 -1515 2140 -1410
rect 3200 -1455 3240 -1400
rect 4250 -930 4290 -920
rect 4250 -1400 4260 -930
rect 4280 -1400 4290 -930
rect 4250 -1410 4290 -1400
rect 5300 -930 5440 -920
rect 5300 -1400 5310 -930
rect 5330 -1400 5360 -930
rect 5380 -1400 5410 -930
rect 5430 -1400 5440 -930
rect 5300 -1410 5440 -1400
rect 6450 -930 6490 -920
rect 6450 -1400 6460 -930
rect 6480 -1400 6490 -930
rect 2195 -1465 3240 -1455
rect 2195 -1485 2205 -1465
rect 2225 -1485 3240 -1465
rect 2195 -1495 3240 -1485
rect 5350 -1515 5390 -1410
rect 2100 -1525 6395 -1515
rect 2100 -1545 6365 -1525
rect 6385 -1545 6395 -1525
rect 2100 -1555 6395 -1545
rect 1000 -1610 2045 -1600
rect 1000 -1630 2015 -1610
rect 2035 -1630 2045 -1610
rect 1000 -1640 2045 -1630
rect -180 -1675 2045 -1665
rect -180 -1695 2015 -1675
rect 2035 -1695 2045 -1675
rect -180 -1705 2045 -1695
rect 2100 -2305 2140 -1555
rect 6450 -1575 6490 -1400
rect 7500 -930 7540 -920
rect 7500 -1400 7510 -930
rect 7530 -1400 7540 -930
rect 7500 -1515 7540 -1400
rect 8550 -930 8690 -920
rect 8550 -1400 8560 -930
rect 8580 -1400 8610 -930
rect 8630 -1400 8660 -930
rect 8680 -1400 8690 -930
rect 8550 -1410 8690 -1400
rect 9700 -930 9740 -920
rect 9700 -1400 9710 -930
rect 9730 -1400 9740 -930
rect 9700 -1410 9740 -1400
rect 10750 -930 10790 -920
rect 10750 -1400 10760 -930
rect 10780 -1400 10790 -930
rect 8605 -1430 8635 -1410
rect 8600 -1440 8640 -1430
rect 8600 -1460 8610 -1440
rect 8630 -1460 8640 -1440
rect 8600 -1470 8640 -1460
rect 6545 -1525 7540 -1515
rect 6545 -1545 6555 -1525
rect 6575 -1545 7540 -1525
rect 6545 -1555 7540 -1545
rect 6450 -1585 8575 -1575
rect 2195 -1610 6395 -1600
rect 2195 -1630 2205 -1610
rect 2225 -1630 6395 -1610
rect 6450 -1605 8545 -1585
rect 8565 -1605 8575 -1585
rect 6450 -1615 8575 -1605
rect 2195 -1640 6395 -1630
rect 6355 -1665 6395 -1640
rect 2195 -1675 5340 -1665
rect 2195 -1695 2205 -1675
rect 2225 -1695 5340 -1675
rect 2195 -1705 5340 -1695
rect 6355 -1705 7540 -1665
rect 3200 -1770 3240 -1750
rect 3150 -1780 3240 -1770
rect 3150 -2250 3160 -1780
rect 3180 -2250 3210 -1780
rect 3230 -2250 3240 -1780
rect 3150 -2260 3240 -2250
rect 4250 -1780 4290 -1770
rect 4250 -2250 4260 -1780
rect 4280 -2250 4290 -1780
rect 4250 -2260 4290 -2250
rect 5300 -1780 5340 -1705
rect 5300 -2250 5310 -1780
rect 5330 -2250 5340 -1780
rect 5300 -2260 5340 -2250
rect 6350 -1780 6490 -1770
rect 6350 -2250 6360 -1780
rect 6380 -2250 6410 -1780
rect 6430 -2250 6460 -1780
rect 6480 -2250 6490 -1780
rect 6350 -2260 6490 -2250
rect 7500 -1780 7540 -1705
rect 8605 -1770 8635 -1470
rect 10750 -1575 10790 -1400
rect 11800 -930 11940 -920
rect 11800 -1400 11810 -930
rect 11830 -1400 11860 -930
rect 11880 -1400 11910 -930
rect 11930 -1400 11940 -930
rect 11800 -1410 11940 -1400
rect 12950 -930 12990 -920
rect 12950 -1400 12960 -930
rect 12980 -1400 12990 -930
rect 11850 -1490 11890 -1410
rect 11850 -1500 12915 -1490
rect 11850 -1520 12885 -1500
rect 12905 -1520 12915 -1500
rect 11850 -1530 12915 -1520
rect 12950 -1575 12990 -1400
rect 14000 -930 14140 -920
rect 14000 -1400 14010 -930
rect 14030 -1400 14060 -930
rect 14080 -1400 14110 -930
rect 14130 -1400 14140 -930
rect 14000 -1410 14140 -1400
rect 15150 -930 15190 -920
rect 15150 -1400 15160 -930
rect 15180 -1400 15190 -930
rect 14050 -1440 14090 -1410
rect 14050 -1460 14060 -1440
rect 14080 -1460 14090 -1440
rect 14050 -1470 14090 -1460
rect 15150 -1490 15190 -1400
rect 16200 -930 16340 -920
rect 16200 -1400 16210 -930
rect 16230 -1400 16260 -930
rect 16280 -1400 16310 -930
rect 16330 -1400 16340 -930
rect 16200 -1410 16340 -1400
rect 17350 -930 17390 -920
rect 17350 -1400 17360 -930
rect 17380 -1400 17390 -930
rect 17350 -1410 17390 -1400
rect 18400 -930 18490 -920
rect 18400 -1400 18410 -930
rect 18430 -1400 18460 -930
rect 18480 -1400 18490 -930
rect 18400 -1410 18490 -1400
rect 13025 -1500 15310 -1490
rect 13025 -1520 13035 -1500
rect 13055 -1520 15310 -1500
rect 13025 -1530 15310 -1520
rect 18550 -1550 18590 -680
rect 8665 -1585 12990 -1575
rect 8665 -1605 8675 -1585
rect 8695 -1605 12990 -1585
rect 8665 -1615 12990 -1605
rect 7500 -2250 7510 -1780
rect 7530 -2250 7540 -1780
rect 7500 -2260 7540 -2250
rect 8550 -1780 8690 -1770
rect 8550 -2250 8560 -1780
rect 8580 -2250 8610 -1780
rect 8630 -2250 8660 -1780
rect 8680 -2250 8690 -1780
rect 8550 -2260 8690 -2250
rect 9700 -1780 9740 -1770
rect 9700 -2250 9710 -1780
rect 9730 -2250 9740 -1780
rect 9700 -2260 9740 -2250
rect 10750 -1780 10890 -1770
rect 10750 -2250 10760 -1780
rect 10780 -2250 10810 -1780
rect 10830 -2250 10860 -1780
rect 10880 -2250 10890 -1780
rect 10750 -2260 10890 -2250
rect 11900 -1780 11940 -1750
rect 11900 -2250 11910 -1780
rect 11930 -2250 11940 -1780
rect 11900 -2260 11940 -2250
rect 12950 -1780 12990 -1770
rect 12950 -2250 12960 -1780
rect 12980 -2250 12990 -1780
rect 8605 -2280 8635 -2260
rect 8600 -2290 8640 -2280
rect 12950 -2290 12990 -2250
rect 14000 -1780 14090 -1770
rect 14000 -2250 14010 -1780
rect 14030 -2250 14060 -1780
rect 14080 -2250 14090 -1780
rect 14000 -2260 14090 -2250
rect 14000 -2280 14040 -2260
rect 2100 -2345 7540 -2305
rect 8600 -2310 8610 -2290
rect 8630 -2310 8640 -2290
rect 8600 -2320 8640 -2310
rect 3200 -2470 3240 -2450
rect 3150 -2480 3240 -2470
rect 3150 -2950 3160 -2480
rect 3180 -2950 3210 -2480
rect 3230 -2950 3240 -2480
rect 3150 -2960 3240 -2950
rect 4250 -2480 4290 -2470
rect 4250 -2950 4260 -2480
rect 4280 -2950 4290 -2480
rect 4250 -2960 4290 -2950
rect 5300 -2480 5340 -2445
rect 5300 -2950 5310 -2480
rect 5330 -2950 5340 -2480
rect 5300 -2960 5340 -2950
rect 6350 -2480 6490 -2470
rect 6350 -2950 6360 -2480
rect 6380 -2950 6410 -2480
rect 6430 -2950 6460 -2480
rect 6480 -2950 6490 -2480
rect 6350 -2960 6490 -2950
rect 7500 -2480 7540 -2345
rect 8605 -2470 8635 -2320
rect 7500 -2950 7510 -2480
rect 7530 -2950 7540 -2480
rect 7500 -2960 7540 -2950
rect 8550 -2480 8690 -2470
rect 8550 -2950 8560 -2480
rect 8580 -2950 8610 -2480
rect 8630 -2950 8660 -2480
rect 8680 -2950 8690 -2480
rect 8550 -2960 8690 -2950
rect 9700 -2480 9740 -2470
rect 9700 -2950 9710 -2480
rect 9730 -2950 9740 -2480
rect 9700 -2960 9740 -2950
rect 10750 -2480 10890 -2470
rect 10750 -2950 10760 -2480
rect 10780 -2950 10810 -2480
rect 10830 -2950 10860 -2480
rect 10880 -2950 10890 -2480
rect 10750 -2960 10890 -2950
rect 11900 -2480 11940 -2450
rect 11900 -2950 11910 -2480
rect 11930 -2950 11940 -2480
rect 11900 -2960 11940 -2950
rect 12950 -2480 12990 -2470
rect 12950 -2950 12960 -2480
rect 12980 -2950 12990 -2480
rect 8605 -2980 8635 -2960
rect 8600 -2990 8640 -2980
rect 12950 -2990 12990 -2950
rect 14000 -2480 14090 -2470
rect 14000 -2950 14010 -2480
rect 14030 -2950 14060 -2480
rect 14080 -2950 14090 -2480
rect 14000 -2960 14090 -2950
rect 14000 -2980 14040 -2960
rect 8600 -3010 8610 -2990
rect 8630 -3010 8640 -2990
rect 8600 -3020 8640 -3010
<< viali >>
rect 6460 -585 6480 -115
rect 12960 -585 12980 -115
rect 4260 -1400 4280 -930
rect 9710 -1400 9730 -930
rect 6360 -2250 6380 -1780
rect 6410 -2250 6430 -1780
rect 6460 -2250 6480 -1780
rect 10760 -2250 10780 -1780
rect 10810 -2250 10830 -1780
rect 10860 -2250 10880 -1780
rect 6360 -2950 6380 -2480
rect 6410 -2950 6430 -2480
rect 6460 -2950 6480 -2480
rect 8560 -2950 8580 -2480
rect 8610 -2950 8630 -2480
rect 8660 -2950 8680 -2480
rect 10760 -2950 10780 -2480
rect 10810 -2950 10830 -2480
rect 10860 -2950 10880 -2480
<< end >>
